// core.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module core (
		input  wire       clk_clk,                          //                       clk.clk
		input  wire       clk_0_clk,                        //                     clk_0.clk
		output wire [9:0] pio_0_external_connection_export, // pio_0_external_connection.export
		input  wire [9:0] pio_1_external_connection_export, // pio_1_external_connection.export
		input  wire       reset_reset_n,                    //                     reset.reset_n
		input  wire       reset_0_reset_n                   //                   reset_0.reset_n
	);

	wire         altpll_0_c0_clk;                                               // altpll_0:c0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, mm_clock_crossing_bridge_1:s0_clk, mm_interconnect_0:altpll_0_c0_clk, mm_interconnect_1:altpll_0_c0_clk, modular_adc_0:adc_pll_clock_clk, nios2_gen2_0:clk, onchip_flash_0:clock, onchip_memory2_0:clk, pio_0:clk, rst_controller_004:clk, timer_0:clk]
	wire         altpll_0_c2_clk;                                               // altpll_0:c2 -> [irq_synchronizer:receiver_clk, mm_clock_crossing_bridge_1:m0_clk, mm_interconnect_1:altpll_0_c2_clk, pio_1:clk, rst_controller_003:clk, sysid_qsys_0:clock]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                             // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                          // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                          // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [24:0] nios2_gen2_0_data_master_address;                              // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                           // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                 // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                        // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                            // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                      // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [24:0] nios2_gen2_0_instruction_master_address;                       // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                          // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_readdata;                 // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	wire   [0:0] mm_interconnect_0_onchip_flash_0_csr_address;                  // mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_0_onchip_flash_0_csr_read;                     // mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire         mm_interconnect_0_onchip_flash_0_csr_write;                    // mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_writedata;                // mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;                // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;             // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire  [18:0] mm_interconnect_0_onchip_flash_0_data_address;                 // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_read;                    // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;           // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_onchip_flash_0_data_write;                   // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;               // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;              // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;       // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;    // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata;      // mm_clock_crossing_bridge_1:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest;   // mm_clock_crossing_bridge_1:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_debugaccess -> mm_clock_crossing_bridge_1:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_address -> mm_clock_crossing_bridge_1:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_read -> mm_clock_crossing_bridge_1:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_byteenable -> mm_clock_crossing_bridge_1:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid; // mm_clock_crossing_bridge_1:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_write -> mm_clock_crossing_bridge_1:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_writedata -> mm_clock_crossing_bridge_1:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_burstcount -> mm_clock_crossing_bridge_1:s0_burstcount
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;              // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                 // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;              // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                   // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;               // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                   // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_modular_adc_0_sample_store_csr_readdata;     // modular_adc_0:sample_store_csr_readdata -> mm_interconnect_0:modular_adc_0_sample_store_csr_readdata
	wire   [6:0] mm_interconnect_0_modular_adc_0_sample_store_csr_address;      // mm_interconnect_0:modular_adc_0_sample_store_csr_address -> modular_adc_0:sample_store_csr_address
	wire         mm_interconnect_0_modular_adc_0_sample_store_csr_read;         // mm_interconnect_0:modular_adc_0_sample_store_csr_read -> modular_adc_0:sample_store_csr_read
	wire         mm_interconnect_0_modular_adc_0_sample_store_csr_write;        // mm_interconnect_0:modular_adc_0_sample_store_csr_write -> modular_adc_0:sample_store_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_0_sample_store_csr_writedata;    // mm_interconnect_0:modular_adc_0_sample_store_csr_writedata -> modular_adc_0:sample_store_csr_writedata
	wire  [31:0] mm_interconnect_0_modular_adc_0_sequencer_csr_readdata;        // modular_adc_0:sequencer_csr_readdata -> mm_interconnect_0:modular_adc_0_sequencer_csr_readdata
	wire   [0:0] mm_interconnect_0_modular_adc_0_sequencer_csr_address;         // mm_interconnect_0:modular_adc_0_sequencer_csr_address -> modular_adc_0:sequencer_csr_address
	wire         mm_interconnect_0_modular_adc_0_sequencer_csr_read;            // mm_interconnect_0:modular_adc_0_sequencer_csr_read -> modular_adc_0:sequencer_csr_read
	wire         mm_interconnect_0_modular_adc_0_sequencer_csr_write;           // mm_interconnect_0:modular_adc_0_sequencer_csr_write -> modular_adc_0:sequencer_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_0_sequencer_csr_writedata;       // mm_interconnect_0:modular_adc_0_sequencer_csr_writedata -> modular_adc_0:sequencer_csr_writedata
	wire         mm_clock_crossing_bridge_1_m0_waitrequest;                     // mm_interconnect_1:mm_clock_crossing_bridge_1_m0_waitrequest -> mm_clock_crossing_bridge_1:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_1_m0_readdata;                        // mm_interconnect_1:mm_clock_crossing_bridge_1_m0_readdata -> mm_clock_crossing_bridge_1:m0_readdata
	wire         mm_clock_crossing_bridge_1_m0_debugaccess;                     // mm_clock_crossing_bridge_1:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_debugaccess
	wire   [9:0] mm_clock_crossing_bridge_1_m0_address;                         // mm_clock_crossing_bridge_1:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_address
	wire         mm_clock_crossing_bridge_1_m0_read;                            // mm_clock_crossing_bridge_1:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_read
	wire   [3:0] mm_clock_crossing_bridge_1_m0_byteenable;                      // mm_clock_crossing_bridge_1:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_byteenable
	wire         mm_clock_crossing_bridge_1_m0_readdatavalid;                   // mm_interconnect_1:mm_clock_crossing_bridge_1_m0_readdatavalid -> mm_clock_crossing_bridge_1:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_1_m0_writedata;                       // mm_clock_crossing_bridge_1:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_writedata
	wire         mm_clock_crossing_bridge_1_m0_write;                           // mm_clock_crossing_bridge_1:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_write
	wire   [0:0] mm_clock_crossing_bridge_1_m0_burstcount;                      // mm_clock_crossing_bridge_1:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_1_m0_burstcount
	wire  [31:0] mm_interconnect_1_sysid_qsys_0_control_slave_readdata;         // sysid_qsys_0:readdata -> mm_interconnect_1:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_qsys_0_control_slave_address;          // mm_interconnect_1:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire         mm_interconnect_1_pio_0_s1_chipselect;                         // mm_interconnect_1:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_1_pio_0_s1_readdata;                           // pio_0:readdata -> mm_interconnect_1:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_0_s1_address;                            // mm_interconnect_1:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_1_pio_0_s1_write;                              // mm_interconnect_1:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_1_pio_0_s1_writedata;                          // mm_interconnect_1:pio_0_s1_writedata -> pio_0:writedata
	wire         mm_interconnect_1_pio_1_s1_chipselect;                         // mm_interconnect_1:pio_1_s1_chipselect -> pio_1:chipselect
	wire  [31:0] mm_interconnect_1_pio_1_s1_readdata;                           // pio_1:readdata -> mm_interconnect_1:pio_1_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_1_s1_address;                            // mm_interconnect_1:pio_1_s1_address -> pio_1:address
	wire         mm_interconnect_1_pio_1_s1_write;                              // mm_interconnect_1:pio_1_s1_write -> pio_1:write_n
	wire  [31:0] mm_interconnect_1_pio_1_s1_writedata;                          // mm_interconnect_1:pio_1_s1_writedata -> pio_1:writedata
	wire         mm_interconnect_1_timer_0_s1_chipselect;                       // mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_1_timer_0_s1_readdata;                         // timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_0_s1_address;                          // mm_interconnect_1:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_1_timer_0_s1_write;                            // mm_interconnect_1:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_1_timer_0_s1_writedata;                        // mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver1_irq;                                      // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                          // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver0_irq;                                      // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                 // pio_1:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> altpll_0:reset
	wire         nios2_gen2_0_debug_reset_request_reset;                        // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2, rst_controller_003:reset_in2, rst_controller_004:reset_in2]
	wire         master_0_master_reset_reset;                                   // master_0:master_reset_reset -> [rst_controller:reset_in3, rst_controller_001:reset_in3, rst_controller_002:reset_in3, rst_controller_003:reset_in3, rst_controller_004:reset_in3]
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [altpll_1:reset, mm_interconnect_0:modular_adc_0_reset_sink_reset_bridge_in_reset_reset, modular_adc_0:reset_sink_reset_n]
	wire         rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> master_0:clk_reset_reset
	wire         rst_controller_003_reset_out_reset;                            // rst_controller_003:reset_out -> [irq_synchronizer:receiver_reset, mm_clock_crossing_bridge_1:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset_reset, pio_1:reset_n, sysid_qsys_0:reset_n]
	wire         rst_controller_004_reset_out_reset;                            // rst_controller_004:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, mm_clock_crossing_bridge_1:s0_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pio_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_flash_0:reset_n, onchip_memory2_0:reset, pio_0:reset_n, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_004_reset_out_reset_req;                        // rst_controller_004:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	core_altpll_0 altpll_0 (
		.clk                (clk_clk),                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (altpll_0_c0_clk),                //                    c0.clk
		.c1                 (),                               //                    c1.clk
		.c2                 (altpll_0_c2_clk),                //                    c2.clk
		.areset             (),                               //        areset_conduit.export
		.locked             (),                               //        locked_conduit.export
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.c3                 (),                               //           (terminated)
		.c4                 (),                               //           (terminated)
		.phasedone          (),                               //           (terminated)
		.phasecounterselect (3'b000),                         //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0)                            //           (terminated)
	);

	core_altpll_1 altpll_1 (
		.clk                (clk_0_clk),                          //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                                   //             pll_slave.read
		.write              (),                                   //                      .write
		.address            (),                                   //                      .address
		.readdata           (),                                   //                      .readdata
		.writedata          (),                                   //                      .writedata
		.c0                 (),                                   //                    c0.clk
		.areset             (),                                   //        areset_conduit.export
		.locked             (),                                   //        locked_conduit.export
		.scandone           (),                                   //           (terminated)
		.scandataout        (),                                   //           (terminated)
		.c1                 (),                                   //           (terminated)
		.c2                 (),                                   //           (terminated)
		.c3                 (),                                   //           (terminated)
		.c4                 (),                                   //           (terminated)
		.phasedone          (),                                   //           (terminated)
		.phasecounterselect (3'b000),                             //           (terminated)
		.phaseupdown        (1'b0),                               //           (terminated)
		.phasestep          (1'b0),                               //           (terminated)
		.scanclk            (1'b0),                               //           (terminated)
		.scanclkena         (1'b0),                               //           (terminated)
		.scandata           (1'b0),                               //           (terminated)
		.configupdate       (1'b0)                                //           (terminated)
	);

	core_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_0_clk),                          //          clk.clk
		.clk_reset_reset      (rst_controller_002_reset_out_reset), //    clk_reset.reset
		.master_address       (),                                   //       master.address
		.master_readdata      (),                                   //             .readdata
		.master_read          (),                                   //             .read
		.master_write         (),                                   //             .write
		.master_writedata     (),                                   //             .writedata
		.master_waitrequest   (),                                   //             .waitrequest
		.master_readdatavalid (),                                   //             .readdatavalid
		.master_byteenable    (),                                   //             .byteenable
		.master_reset_reset   (master_0_master_reset_reset)         // master_reset.reset
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_1 (
		.m0_clk           (altpll_0_c2_clk),                                               //   m0_clk.clk
		.m0_reset         (rst_controller_003_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (altpll_0_c0_clk),                                               //   s0_clk.clk
		.s0_reset         (rst_controller_004_reset_out_reset),                            // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_1_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_1_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_1_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_1_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_1_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_1_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_1_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_1_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_1_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_1_m0_debugaccess)                      //         .debugaccess
	);

	core_modular_adc_0 #(
		.is_this_first_or_second_adc (1)
	) modular_adc_0 (
		.clock_clk                  (clk_0_clk),                                                  //            clock.clk
		.reset_sink_reset_n         (~rst_controller_001_reset_out_reset),                        //       reset_sink.reset_n
		.adc_pll_clock_clk          (altpll_0_c0_clk),                                            //    adc_pll_clock.clk
		.adc_pll_locked_export      (),                                                           //   adc_pll_locked.export
		.sequencer_csr_address      (mm_interconnect_0_modular_adc_0_sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (mm_interconnect_0_modular_adc_0_sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (mm_interconnect_0_modular_adc_0_sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (mm_interconnect_0_modular_adc_0_sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (mm_interconnect_0_modular_adc_0_sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (mm_interconnect_0_modular_adc_0_sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (mm_interconnect_0_modular_adc_0_sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (mm_interconnect_0_modular_adc_0_sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (mm_interconnect_0_modular_adc_0_sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (mm_interconnect_0_modular_adc_0_sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       ()                                                            // sample_store_irq.irq
	);

	core_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_004_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_004_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M50DAF484C6GES"),
		.DEVICE_ID                           ("50"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (8191),
		.SECTOR2_START_ADDR                  (8192),
		.SECTOR2_END_ADDR                    (16383),
		.SECTOR3_START_ADDR                  (16384),
		.SECTOR3_END_ADDR                    (114687),
		.SECTOR4_START_ADDR                  (114688),
		.SECTOR4_END_ADDR                    (188415),
		.SECTOR5_START_ADDR                  (188416),
		.SECTOR5_END_ADDR                    (360447),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (360447),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (16383),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (360447),
		.ADDR_RANGE2_END_ADDR                (360447),
		.ADDR_RANGE1_OFFSET                  (2048),
		.ADDR_RANGE2_OFFSET                  (0),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (19),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (0),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (5),
		.FLASH_RESET_CYCLE_MAX_INDEX         (20),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (96),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (28000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (24400),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("False"),
		.IS_COMPRESSED_IMAGE                 ("False")
	) onchip_flash_0 (
		.clock                   (altpll_0_c0_clk),                                     //    clk.clk
		.reset_n                 (~rst_controller_004_reset_out_reset),                 // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_onchip_flash_0_csr_readdata)        //       .readdata
	);

	core_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_004_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_004_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	core_pio_0 pio_0 (
		.clk        (altpll_0_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_1_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)       // external_connection.export
	);

	core_pio_1 pio_1 (
		.clk        (altpll_0_c2_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_1_pio_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_1_s1_readdata),   //                    .readdata
		.in_port    (pio_1_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)          //                 irq.irq
	);

	core_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c2_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_0_control_slave_address)   //              .address
	);

	core_timer_0 timer_0 (
		.clk        (altpll_0_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_1_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	core_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                      (altpll_0_c0_clk),                                               //                                    altpll_0_c0.clk
		.clk_1_clk_clk                                        (clk_0_clk),                                                     //                                      clk_1_clk.clk
		.modular_adc_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                            // modular_adc_0_reset_sink_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset       (rst_controller_004_reset_out_reset),                            //       nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                     (nios2_gen2_0_data_master_address),                              //                       nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                 (nios2_gen2_0_data_master_waitrequest),                          //                                               .waitrequest
		.nios2_gen2_0_data_master_byteenable                  (nios2_gen2_0_data_master_byteenable),                           //                                               .byteenable
		.nios2_gen2_0_data_master_read                        (nios2_gen2_0_data_master_read),                                 //                                               .read
		.nios2_gen2_0_data_master_readdata                    (nios2_gen2_0_data_master_readdata),                             //                                               .readdata
		.nios2_gen2_0_data_master_readdatavalid               (nios2_gen2_0_data_master_readdatavalid),                        //                                               .readdatavalid
		.nios2_gen2_0_data_master_write                       (nios2_gen2_0_data_master_write),                                //                                               .write
		.nios2_gen2_0_data_master_writedata                   (nios2_gen2_0_data_master_writedata),                            //                                               .writedata
		.nios2_gen2_0_data_master_debugaccess                 (nios2_gen2_0_data_master_debugaccess),                          //                                               .debugaccess
		.nios2_gen2_0_instruction_master_address              (nios2_gen2_0_instruction_master_address),                       //                nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest          (nios2_gen2_0_instruction_master_waitrequest),                   //                                               .waitrequest
		.nios2_gen2_0_instruction_master_read                 (nios2_gen2_0_instruction_master_read),                          //                                               .read
		.nios2_gen2_0_instruction_master_readdata             (nios2_gen2_0_instruction_master_readdata),                      //                                               .readdata
		.nios2_gen2_0_instruction_master_readdatavalid        (nios2_gen2_0_instruction_master_readdatavalid),                 //                                               .readdatavalid
		.mm_clock_crossing_bridge_1_s0_address                (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address),       //                  mm_clock_crossing_bridge_1_s0.address
		.mm_clock_crossing_bridge_1_s0_write                  (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write),         //                                               .write
		.mm_clock_crossing_bridge_1_s0_read                   (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read),          //                                               .read
		.mm_clock_crossing_bridge_1_s0_readdata               (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata),      //                                               .readdata
		.mm_clock_crossing_bridge_1_s0_writedata              (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata),     //                                               .writedata
		.mm_clock_crossing_bridge_1_s0_burstcount             (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount),    //                                               .burstcount
		.mm_clock_crossing_bridge_1_s0_byteenable             (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable),    //                                               .byteenable
		.mm_clock_crossing_bridge_1_s0_readdatavalid          (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid), //                                               .readdatavalid
		.mm_clock_crossing_bridge_1_s0_waitrequest            (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest),   //                                               .waitrequest
		.mm_clock_crossing_bridge_1_s0_debugaccess            (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess),   //                                               .debugaccess
		.modular_adc_0_sample_store_csr_address               (mm_interconnect_0_modular_adc_0_sample_store_csr_address),      //                 modular_adc_0_sample_store_csr.address
		.modular_adc_0_sample_store_csr_write                 (mm_interconnect_0_modular_adc_0_sample_store_csr_write),        //                                               .write
		.modular_adc_0_sample_store_csr_read                  (mm_interconnect_0_modular_adc_0_sample_store_csr_read),         //                                               .read
		.modular_adc_0_sample_store_csr_readdata              (mm_interconnect_0_modular_adc_0_sample_store_csr_readdata),     //                                               .readdata
		.modular_adc_0_sample_store_csr_writedata             (mm_interconnect_0_modular_adc_0_sample_store_csr_writedata),    //                                               .writedata
		.modular_adc_0_sequencer_csr_address                  (mm_interconnect_0_modular_adc_0_sequencer_csr_address),         //                    modular_adc_0_sequencer_csr.address
		.modular_adc_0_sequencer_csr_write                    (mm_interconnect_0_modular_adc_0_sequencer_csr_write),           //                                               .write
		.modular_adc_0_sequencer_csr_read                     (mm_interconnect_0_modular_adc_0_sequencer_csr_read),            //                                               .read
		.modular_adc_0_sequencer_csr_readdata                 (mm_interconnect_0_modular_adc_0_sequencer_csr_readdata),        //                                               .readdata
		.modular_adc_0_sequencer_csr_writedata                (mm_interconnect_0_modular_adc_0_sequencer_csr_writedata),       //                                               .writedata
		.nios2_gen2_0_debug_mem_slave_address                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),        //                   nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),          //                                               .write
		.nios2_gen2_0_debug_mem_slave_read                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),           //                                               .read
		.nios2_gen2_0_debug_mem_slave_readdata                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),       //                                               .readdata
		.nios2_gen2_0_debug_mem_slave_writedata               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),      //                                               .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),     //                                               .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),    //                                               .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),    //                                               .debugaccess
		.onchip_flash_0_csr_address                           (mm_interconnect_0_onchip_flash_0_csr_address),                  //                             onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                             (mm_interconnect_0_onchip_flash_0_csr_write),                    //                                               .write
		.onchip_flash_0_csr_read                              (mm_interconnect_0_onchip_flash_0_csr_read),                     //                                               .read
		.onchip_flash_0_csr_readdata                          (mm_interconnect_0_onchip_flash_0_csr_readdata),                 //                                               .readdata
		.onchip_flash_0_csr_writedata                         (mm_interconnect_0_onchip_flash_0_csr_writedata),                //                                               .writedata
		.onchip_flash_0_data_address                          (mm_interconnect_0_onchip_flash_0_data_address),                 //                            onchip_flash_0_data.address
		.onchip_flash_0_data_write                            (mm_interconnect_0_onchip_flash_0_data_write),                   //                                               .write
		.onchip_flash_0_data_read                             (mm_interconnect_0_onchip_flash_0_data_read),                    //                                               .read
		.onchip_flash_0_data_readdata                         (mm_interconnect_0_onchip_flash_0_data_readdata),                //                                               .readdata
		.onchip_flash_0_data_writedata                        (mm_interconnect_0_onchip_flash_0_data_writedata),               //                                               .writedata
		.onchip_flash_0_data_burstcount                       (mm_interconnect_0_onchip_flash_0_data_burstcount),              //                                               .burstcount
		.onchip_flash_0_data_readdatavalid                    (mm_interconnect_0_onchip_flash_0_data_readdatavalid),           //                                               .readdatavalid
		.onchip_flash_0_data_waitrequest                      (mm_interconnect_0_onchip_flash_0_data_waitrequest),             //                                               .waitrequest
		.onchip_memory2_0_s1_address                          (mm_interconnect_0_onchip_memory2_0_s1_address),                 //                            onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                            (mm_interconnect_0_onchip_memory2_0_s1_write),                   //                                               .write
		.onchip_memory2_0_s1_readdata                         (mm_interconnect_0_onchip_memory2_0_s1_readdata),                //                                               .readdata
		.onchip_memory2_0_s1_writedata                        (mm_interconnect_0_onchip_memory2_0_s1_writedata),               //                                               .writedata
		.onchip_memory2_0_s1_byteenable                       (mm_interconnect_0_onchip_memory2_0_s1_byteenable),              //                                               .byteenable
		.onchip_memory2_0_s1_chipselect                       (mm_interconnect_0_onchip_memory2_0_s1_chipselect),              //                                               .chipselect
		.onchip_memory2_0_s1_clken                            (mm_interconnect_0_onchip_memory2_0_s1_clken)                    //                                               .clken
	);

	core_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c0_clk                                                 (altpll_0_c0_clk),                                       //                                               altpll_0_c0.clk
		.altpll_0_c2_clk                                                 (altpll_0_c2_clk),                                       //                                               altpll_0_c2.clk
		.mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                    // mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset.reset
		.pio_0_reset_reset_bridge_in_reset_reset                         (rst_controller_004_reset_out_reset),                    //                         pio_0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_1_m0_address                           (mm_clock_crossing_bridge_1_m0_address),                 //                             mm_clock_crossing_bridge_1_m0.address
		.mm_clock_crossing_bridge_1_m0_waitrequest                       (mm_clock_crossing_bridge_1_m0_waitrequest),             //                                                          .waitrequest
		.mm_clock_crossing_bridge_1_m0_burstcount                        (mm_clock_crossing_bridge_1_m0_burstcount),              //                                                          .burstcount
		.mm_clock_crossing_bridge_1_m0_byteenable                        (mm_clock_crossing_bridge_1_m0_byteenable),              //                                                          .byteenable
		.mm_clock_crossing_bridge_1_m0_read                              (mm_clock_crossing_bridge_1_m0_read),                    //                                                          .read
		.mm_clock_crossing_bridge_1_m0_readdata                          (mm_clock_crossing_bridge_1_m0_readdata),                //                                                          .readdata
		.mm_clock_crossing_bridge_1_m0_readdatavalid                     (mm_clock_crossing_bridge_1_m0_readdatavalid),           //                                                          .readdatavalid
		.mm_clock_crossing_bridge_1_m0_write                             (mm_clock_crossing_bridge_1_m0_write),                   //                                                          .write
		.mm_clock_crossing_bridge_1_m0_writedata                         (mm_clock_crossing_bridge_1_m0_writedata),               //                                                          .writedata
		.mm_clock_crossing_bridge_1_m0_debugaccess                       (mm_clock_crossing_bridge_1_m0_debugaccess),             //                                                          .debugaccess
		.pio_0_s1_address                                                (mm_interconnect_1_pio_0_s1_address),                    //                                                  pio_0_s1.address
		.pio_0_s1_write                                                  (mm_interconnect_1_pio_0_s1_write),                      //                                                          .write
		.pio_0_s1_readdata                                               (mm_interconnect_1_pio_0_s1_readdata),                   //                                                          .readdata
		.pio_0_s1_writedata                                              (mm_interconnect_1_pio_0_s1_writedata),                  //                                                          .writedata
		.pio_0_s1_chipselect                                             (mm_interconnect_1_pio_0_s1_chipselect),                 //                                                          .chipselect
		.pio_1_s1_address                                                (mm_interconnect_1_pio_1_s1_address),                    //                                                  pio_1_s1.address
		.pio_1_s1_write                                                  (mm_interconnect_1_pio_1_s1_write),                      //                                                          .write
		.pio_1_s1_readdata                                               (mm_interconnect_1_pio_1_s1_readdata),                   //                                                          .readdata
		.pio_1_s1_writedata                                              (mm_interconnect_1_pio_1_s1_writedata),                  //                                                          .writedata
		.pio_1_s1_chipselect                                             (mm_interconnect_1_pio_1_s1_chipselect),                 //                                                          .chipselect
		.sysid_qsys_0_control_slave_address                              (mm_interconnect_1_sysid_qsys_0_control_slave_address),  //                                sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                             (mm_interconnect_1_sysid_qsys_0_control_slave_readdata), //                                                          .readdata
		.timer_0_s1_address                                              (mm_interconnect_1_timer_0_s1_address),                  //                                                timer_0_s1.address
		.timer_0_s1_write                                                (mm_interconnect_1_timer_0_s1_write),                    //                                                          .write
		.timer_0_s1_readdata                                             (mm_interconnect_1_timer_0_s1_readdata),                 //                                                          .readdata
		.timer_0_s1_writedata                                            (mm_interconnect_1_timer_0_s1_writedata),                //                                                          .writedata
		.timer_0_s1_chipselect                                           (mm_interconnect_1_timer_0_s1_chipselect)                //                                                          .chipselect
	);

	core_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c2_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (~reset_0_reset_n),                       // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_0_reset_n),                       // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (clk_0_clk),                              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_0_reset_n),                       // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (),                                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (~reset_0_reset_n),                       // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (altpll_0_c2_clk),                        //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (~reset_0_reset_n),                       // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
